// Sample Verilog
module example();
    initial begin
        $display("Hello VLSI!");
    end
endmodule
