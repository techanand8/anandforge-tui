// Mayank Design
